* SPICE3 file created from inverter.ext - technology: sky130A

.option scale=10m

Vpower vdd gnd 3.3
Vin A gnd pulse(0, 3.3, 100p, 50p, 200p, 500p)

X0 Vout Vin Gnd Gnd sky130_fd_pr__nfet_01v8 ad=4.75n pd=0.29m as=4.75n ps=0.29m w=95 l=15
X1 Vout Vin Vdd Vdd sky130_fd_pr__pfet_01v8 ad=4.75n pd=0.29m as=4.75n ps=0.29m w=95 l=15

.tran 1p 1200p
.end
