magic
tech scmos
timestamp 1752860621
<< nwell >>
rect -6 -6 48 14
rect 59 -6 96 14
<< ntransistor >>
rect 11 -26 14 -18
rect 28 -26 31 -18
rect 76 -26 79 -18
<< ptransistor >>
rect 11 0 14 8
rect 28 0 31 8
rect 76 0 79 8
<< ndiffusion >>
rect 0 -19 11 -18
rect 0 -25 1 -19
rect 7 -25 11 -19
rect 0 -26 11 -25
rect 14 -26 28 -18
rect 31 -19 42 -18
rect 31 -25 35 -19
rect 41 -25 42 -19
rect 31 -26 42 -25
rect 65 -19 76 -18
rect 65 -25 66 -19
rect 72 -25 76 -19
rect 65 -26 76 -25
rect 79 -19 90 -18
rect 79 -25 83 -19
rect 89 -25 90 -19
rect 79 -26 90 -25
<< pdiffusion >>
rect 0 7 11 8
rect 0 1 1 7
rect 7 1 11 7
rect 0 0 11 1
rect 14 7 28 8
rect 14 1 18 7
rect 24 1 28 7
rect 14 0 28 1
rect 31 7 42 8
rect 31 1 35 7
rect 41 1 42 7
rect 31 0 42 1
rect 65 7 76 8
rect 65 1 66 7
rect 72 1 76 7
rect 65 0 76 1
rect 79 7 90 8
rect 79 1 83 7
rect 89 1 90 7
rect 79 0 90 1
<< ndcontact >>
rect 1 -25 7 -19
rect 35 -25 41 -19
rect 66 -25 72 -19
rect 83 -25 89 -19
<< pdcontact >>
rect 1 1 7 7
rect 18 1 24 7
rect 35 1 41 7
rect 66 1 72 7
rect 83 1 89 7
<< psubstratepcontact >>
rect 18 -38 24 -32
rect 49 -38 55 -32
<< nsubstratencontact >>
rect 18 20 24 26
rect 52 20 58 26
<< polysilicon >>
rect 11 8 14 11
rect 28 8 31 11
rect 76 8 79 11
rect 11 -18 14 0
rect 28 -18 31 0
rect 76 -9 79 0
rect 72 -15 79 -9
rect 76 -18 79 -15
rect 11 -29 14 -26
rect 28 -29 31 -26
rect 76 -29 79 -26
<< polycontact >>
rect 66 -15 72 -9
<< metal1 >>
rect 1 20 18 26
rect 24 20 52 26
rect 58 20 72 26
rect 1 7 7 20
rect 35 7 41 20
rect 66 7 72 20
rect 18 -9 24 1
rect 83 -9 89 1
rect 18 -15 66 -9
rect 83 -15 95 -9
rect 35 -19 41 -15
rect 83 -19 89 -15
rect 1 -32 7 -25
rect 66 -32 72 -25
rect 1 -38 18 -32
rect 24 -38 49 -32
rect 55 -38 72 -32
<< labels >>
rlabel polysilicon 12 -17 12 -17 1 A
rlabel polysilicon 29 -17 29 -17 1 B
rlabel metal1 92 -12 92 -12 7 Z
rlabel metal1 38 23 38 23 5 vdd
rlabel metal1 38 -35 38 -35 1 gnd
<< end >>
