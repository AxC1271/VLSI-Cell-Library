* SPICE3 file created from /home/parallels/Documents/vlsi_layouts/logic_gates/nor_gate/nor_gate.ext - technology: scmos

.include ./ami05.txt
.option scale=0.3u
.options method=gear reltol=1e-4 abstol=1e-12 vabstol=1e-12

* Power
Vdd vdd 0 3.3

* Input Pulses
VA A 0 PULSE(0 3.3 5n 1p 1p 5n 10n)
VB B 0 PULSE(0 3.3 10n 1p 1p 10n 20n)

* NOR Gate

M1000 gnd B Z Gnd nfet w=8 l=3
+  ad=176 pd=76 as=112 ps=44
M1001 Z B a_14_0# w_n6_n6# pfet w=8 l=3
+  ad=88 pd=38 as=112 ps=44
M1002 a_14_0# A vdd w_n6_n6# pfet w=8 l=3
+  ad=0 pd=0 as=88 ps=38
M1003 Z A gnd Gnd nfet w=8 l=3
+  ad=0 pd=0 as=0 ps=0

* Parasitics
C0 0 0 3.47fF
C1 vdd 2.04fF
C2 w_n6_n6# 0 3.89fF
Cload Z 0 80f

.tran 1n 40n

.end
