magic
tech scmos
timestamp 1759099264
<< nwell >>
rect -6 -6 48 14
<< ntransistor >>
rect 11 -22 14 -14
rect 28 -22 31 -14
<< ptransistor >>
rect 11 0 14 8
rect 28 0 31 8
<< ndiffusion >>
rect 0 -15 11 -14
rect 0 -21 1 -15
rect 7 -21 11 -15
rect 0 -22 11 -21
rect 14 -22 28 -14
rect 31 -15 42 -14
rect 31 -21 35 -15
rect 41 -21 42 -15
rect 31 -22 42 -21
<< pdiffusion >>
rect 0 7 11 8
rect 0 1 1 7
rect 7 1 11 7
rect 0 0 11 1
rect 14 7 28 8
rect 14 1 18 7
rect 24 1 28 7
rect 14 0 28 1
rect 31 7 42 8
rect 31 1 35 7
rect 41 1 42 7
rect 31 0 42 1
<< ndcontact >>
rect 1 -21 7 -15
rect 35 -21 41 -15
<< pdcontact >>
rect 1 1 7 7
rect 18 1 24 7
rect 35 1 41 7
<< psubstratepcontact >>
rect 18 -39 24 -33
<< nsubstratencontact >>
rect 18 22 24 28
<< polysilicon >>
rect 11 8 14 11
rect 28 8 31 11
rect 11 -14 14 0
rect 28 -14 31 0
rect 11 -25 14 -22
rect 28 -25 31 -22
<< metal1 >>
rect 1 22 18 28
rect 24 22 41 28
rect 1 7 7 22
rect 35 7 41 22
rect 18 -7 24 1
rect 18 -12 47 -7
rect 35 -15 41 -12
rect 1 -33 7 -21
rect 1 -39 18 -33
rect 24 -39 31 -33
<< labels >>
rlabel metal1 15 -36 15 -36 1 gnd
rlabel metal1 15 25 15 25 5 vdd
rlabel polysilicon 12 -13 12 -13 1 A
rlabel polysilicon 29 -13 29 -13 1 B
rlabel metal1 44 -10 44 -10 7 Z
<< end >>
