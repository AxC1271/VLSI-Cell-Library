magic
tech scmos
timestamp 1759165093
<< polysilicon >>
rect 44 4 47 9
rect 110 4 113 9
rect 44 -71 47 -66
rect 110 -71 113 -66
<< polycontact >>
rect 22 22 27 27
rect 88 22 93 27
rect 47 4 53 10
rect 113 4 118 9
rect 22 -53 27 -48
rect 88 -53 93 -48
rect 47 -71 52 -66
rect 113 -71 118 -66
<< metal1 >>
rect 63 22 88 27
rect 129 22 150 27
rect 53 9 59 10
rect 53 5 54 9
rect 58 5 59 9
rect 53 4 59 5
rect 0 -7 14 -6
rect 0 -11 9 -7
rect 13 -11 14 -7
rect 0 -12 14 -11
rect 0 -48 5 -12
rect 67 -39 73 22
rect 118 4 140 9
rect 67 -43 68 -39
rect 72 -43 73 -39
rect 67 -44 73 -43
rect 135 -48 140 4
rect 0 -53 22 -48
rect 63 -53 88 -48
rect 129 -53 140 -48
rect 67 -58 73 -57
rect 67 -62 68 -58
rect 72 -62 73 -58
rect 67 -66 73 -62
rect 145 -66 150 22
rect 52 -71 73 -66
rect 118 -71 150 -66
<< m2contact >>
rect 54 5 58 9
rect 9 -11 13 -7
rect 68 -43 72 -39
rect 68 -62 72 -58
<< metal2 >>
rect 53 9 59 10
rect 53 5 54 9
rect 58 5 59 9
rect 53 -6 59 5
rect 8 -7 59 -6
rect 8 -11 9 -7
rect 13 -11 59 -7
rect 8 -12 59 -11
rect 67 -39 73 -38
rect 67 -43 68 -39
rect 72 -43 73 -39
rect 67 -58 73 -43
rect 67 -62 68 -58
rect 72 -62 73 -58
rect 67 -63 73 -62
use nand_gate  nand_gate_0 ~/Documents/vlsi_layouts/logic_gates/nand_gate
timestamp 1759099264
transform 1 0 16 0 1 34
box -6 -39 48 28
use nand_gate  nand_gate_1
timestamp 1759099264
transform 1 0 16 0 1 -41
box -6 -39 48 28
use nand_gate  nand_gate_2
timestamp 1759099264
transform 1 0 82 0 1 34
box -6 -39 48 28
use nand_gate  nand_gate_3
timestamp 1759099264
transform 1 0 82 0 1 -41
box -6 -39 48 28
<< labels >>
rlabel polycontact 51 8 51 8 1 en
rlabel polycontact 24 24 24 24 1 d
rlabel metal1 148 25 148 25 7 Q
rlabel metal1 138 -51 138 -51 1 Q_not
<< end >>
