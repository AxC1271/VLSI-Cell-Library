* SPICE3 file created from /home/parallels/Documents/vlsi_layouts/logic_gates/or_gate/or_gate.ext - technology: scmos

.include ./ami05.txt
.option scale=0.3u
.options method=gear reltol=1e-4 abstol=1e-12 vabstol=1e-12

* Power
Vdd vdd 0 3.3

* Input Pulses
VA A 0 PULSE(0 3.3 5n 1p 1p 5n 10n)
VB B 0 PULSE(0 3.3 10n 1p 1p 10n 20n)

* OR Gate
M1000 gnd B a_14_n26# Gnd nfet w=8 l=3
+  ad=264 pd=114 as=112 ps=44
M1001 a_14_n26# B a_14_0# w_n6_n6# pfet w=8 l=3
+  ad=88 pd=38 as=112 ps=44
M1002 Z a_14_n26# vdd w_58_n6# pfet w=8 l=3
+  ad=88 pd=38 as=176 ps=76
M1003 a_14_0# A vdd w_n6_n6# pfet w=8 l=3
+  ad=0 pd=0 as=0 ps=0
M1004 a_14_n26# A gnd Gnd nfet w=8 l=3
+  ad=0 pd=0 as=0 ps=0
M1005 Z a_14_n26# gnd Gnd nfet w=8 l=3
+  ad=88 pd=38 as=0 ps=0

* Parasitics
C0 gnd Gnd 4.75fF
C1 a_14_n26# Gnd 3.79fF
C2 vdd Gnd 4.53fF
C3 w_58_n6# Gnd 2.38fF
C4 w_n6_n6# Gnd 3.89fF

.tran 1n 40n
.end
